module debounce (q,u,n,b,d,led1,led2);
		input wire q,u,n,b,           //四位开关作为密码输入
		input wire d,				  //一位按键作为开锁使能信号
		output wire led1,    	      //保险箱打开信号对应的led输出
		output wire led2			  //报警信号对应的led输出
	wire  [3:0]   code;			  //四位变量存储密码
	reg			  open;			  //保险箱开箱信号
	reg			  alarm;          //报警信号
	assign		code = {q,u,n,b};
	always@(d or code)
		if(d == 1'b1)             //使能，开始判断密码
			begin
				if(code == 4'b0101)   
					begin
					open = 1'b1;  //开锁
					alarm = 1'b0; //没报警
					end
				else
					begin
					open = 1'b0;  
					alarm = 1'b1;
					end
			end
		else
			begin
			open = 1'b0;
			end
	assign  led1 = ~open;		//led亮表示密码锁没开
	assign	led2 = ~alarm;		//led亮代表发出报警信号
endmodule
